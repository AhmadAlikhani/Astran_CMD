.SUBCKT XNOR3 A B C OUT GND VCC
M0P OUT ^C VCC VCC pmos L=65n W=800n 
M1N GND ^C OUT GND nmos L=65n W=480n
.ENDS XNOR3 
