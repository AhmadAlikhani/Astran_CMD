magic
tech scmos
magscale 1 2
timestamp 1687299807
<< m2contact >>
rect 164 674 198 708
<< m2contact >>
rect 164 600 198 634
<< m2contact >>
rect 172 304 206 338
<< m2contact >>
rect 128 434 162 468
<< m2contact >>
rect 64 674 98 708
<< m2contact >>
rect 64 600 98 634
<< m2contact >>
rect 72 304 106 338
<< poly >>
rect 120 464 144 488
<< poly >>
rect 118 464 144 776
<< poly >>
rect 126 414 150 438
<< poly >>
rect 120 414 170 488
<< poly >>
rect 126 412 150 436
<< poly >>
rect 126 412 150 438
<< poly >>
rect 126 236 152 436
<< ndiff >>
rect 168 288 210 384
<< ndiff >>
rect 68 288 210 384
<< ndiff >>
rect 68 288 110 384
<< pdiff >>
rect 160 516 202 724
<< pdiff >>
rect 60 516 202 724
<< pdiff >>
rect 60 516 102 724
<< ndiffusion >>
rect -36 -36 276 456
<< pdiffusion >>
rect -36 456 276 1076
<< nwell >>
rect -94 456 334 1134
<< pwell >>
rect -94 -94 334 456
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 936
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 588 202 720
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 292 208 350
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 104 208 332
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 128 416 206 500
<< metal1 >>
rect 44 300 84 640
<< metal1 >>
rect 44 600 110 708
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 60 300 100 340
<< metal1 >>
rect 44 300 112 340
<< metal1 >>
rect 60 300 118 340
<< glass >>
rect 0 0 240 1040
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 60 300 118 340
<< metal1 >>
rect 44 300 112 340
<< metal1 >>
rect 60 300 100 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 600 110 708
<< metal1 >>
rect 44 300 84 640
<< metal1 >>
rect 128 416 206 500
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 104 208 332
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 168 292 208 350
<< metal1 >>
rect 168 292 208 332
<< metal1 >>
rect 162 588 202 720
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 162 680 202 936
<< metal1 >>
rect 162 680 202 720
<< metal1 >>
rect 140 460 180 500
<< metal1 >>
rect 60 300 100 340
<< end >>