magic
tech scmos
timestamp 1684523853
<< m2contact >>
rect -2 -2 2 2
<< end >>
