magic
tech scmos
magscale 1 2
timestamp 1686780763
<< m2contact >>
rect 164 674 198 708
<< m2contact >>
rect 164 600 198 634
<< m2contact >>
rect 160 304 194 338
<< m2contact >>
rect 128 434 162 468
<< m2contact >>
rect 64 674 98 708
<< m2contact >>
rect 64 600 98 634
<< m2contact >>
rect 60 304 94 338
<< poly >>
rect 120 464 144 488
<< poly >>
rect 118 464 144 776
<< poly >>
rect 120 412 144 436
<< poly >>
rect 120 412 170 488
<< poly >>
rect 116 412 140 436
<< poly >>
rect 116 412 144 436
<< poly >>
rect 114 236 140 436
<< ndiff >>
rect 156 288 198 384
<< ndiff >>
rect 56 288 198 384
<< ndiff >>
rect 56 288 98 384
<< pdiff >>
rect 160 516 202 724
<< pdiff >>
rect 60 516 202 724
<< pdiff >>
rect 60 516 102 724
<< ndiffusion >>
rect -36 -36 276 456
<< pdiffusion >>
rect -36 456 276 1076
<< nwell >>
rect -94 456 334 1134
<< pwell >>
rect -94 -94 334 456
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 936
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 588 204 720
<< metal1 >>
rect 160 104 200 332
<< metal1 >>
rect 160 292 200 350
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 128 416 206 500
<< metal1 >>
rect 44 300 84 640
<< metal1 >>
rect 44 600 110 708
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 66 300 106 340
<< metal1 >>
rect 44 300 112 340
<< metal1 >>
rect 48 300 106 340
<< glass >>
rect 0 0 240 1040
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 48 300 106 340
<< metal1 >>
rect 44 300 112 340
<< metal1 >>
rect 66 300 106 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 300 84 340
<< metal1 >>
rect 44 600 110 708
<< metal1 >>
rect 44 300 84 640
<< metal1 >>
rect 128 416 206 500
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 292 200 350
<< metal1 >>
rect 160 104 200 332
<< metal1 >>
rect 164 588 204 720
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 936
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 140 460 180 500
<< metal1 >>
rect 60 300 100 340
<< end >>