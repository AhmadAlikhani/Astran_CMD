magic
tech scmos
timestamp 1684523853
<< end >>
