magic
tech scmos
magscale 1 2
timestamp 1684523853
<< ndiffusion >>
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
<< end >>
