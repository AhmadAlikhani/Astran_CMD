.SUBCKT XNOR2_CMOS A Q GND VCC
MN Q A GND GND nmos L=65n W=480n
MP Q A VCC VCC pmos L=65n W=800n
.ENDS XNOR2_CMOS 
