magic
tech scmos
magscale 1 2
timestamp 1686778612
<< contact >>
rect 160 572 194 606
<< contact >>
rect 160 306 194 340
<< contact >>
rect 132 436 166 470
<< contact >>
rect 60 572 94 606
<< contact >>
rect 60 306 94 340
<< poly >>
rect 116 466 140 490
<< poly >>
rect 114 466 140 674
<< poly >>
rect 116 416 140 440
<< poly >>
rect 116 416 174 490
<< poly >>
rect 116 384 140 440
<< poly >>
rect 116 416 140 440
<< poly >>
rect 114 250 140 408
<< ndiff >>
rect 144 302 210 356
<< ndiff >>
rect 44 302 210 356
<< ndiff >>
rect 44 302 110 356
<< pdiff >>
rect 156 518 198 622
<< pdiff >>
rect 56 518 198 622
<< pdiff >>
rect 56 518 98 622
<< ndiffusion >>
rect -36 -36 276 456
<< pdiffusion >>
rect -36 456 276 1076
<< nwell >>
rect -94 456 334 1134
<< pwell >>
rect -94 -94 334 456
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 578 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 560 200 618
<< metal1 >>
rect 160 104 200 334
<< metal1 >>
rect 160 294 200 352
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 132 424 208 512
<< metal1 >>
rect 48 300 88 606
<< metal1 >>
rect 48 566 106 606
<< metal1 >>
rect 48 300 88 340
<< metal1 >>
rect 48 300 88 340
<< metal1 >>
rect 54 300 94 340
<< metal1 >>
rect 48 300 112 340
<< metal1 >>
rect 48 300 106 340
<< glass >>
rect 0 0 240 1040
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 48 300 106 340
<< metal1 >>
rect 48 300 112 340
<< metal1 >>
rect 54 300 94 340
<< metal1 >>
rect 48 300 88 340
<< metal1 >>
rect 48 300 88 340
<< metal1 >>
rect 48 566 106 606
<< metal1 >>
rect 48 300 88 606
<< metal1 >>
rect 132 424 208 512
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 104 200 144
<< metal1 >>
rect 160 294 200 352
<< metal1 >>
rect 160 104 200 334
<< metal1 >>
rect 160 560 200 618
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 578 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 160 896 200 936
<< metal1 >>
rect 140 460 180 500
<< metal1 >>
rect 60 300 100 340
<< end >>