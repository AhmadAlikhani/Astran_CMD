magic
tech scmos
magscale 1 2
timestamp 1684523853
<< m2contact >>
<< genericcontact >>
rect 164 674 198 708
<< poly >>
rect 164 600 198 634
<< pdiff >>
rect 160 304 194 338
<< ndiffusion >>
rect 128 434 162 468
<< pdiffusion >>
rect 64 674 98 708
<< nwell >>
rect 64 600 98 634
<< via >>
rect 60 304 94 338
<< genericcontact >>
rect 120 464 144 488
<< poly >>
rect 118 464 144 776
<< ndiff >>
rect 120 412 144 436
<< pdiff >>
rect 120 412 170 488
<< ndiffusion >>
rect 116 412 140 436
<< pdiffusion >>
rect 116 412 144 436
<< nwell >>
rect 114 236 140 436
<< genericcontact >>
rect 156 288 198 384
<< poly >>
rect 56 288 198 384
<< ndiff >>
rect 56 288 98 384
<< genericcontact >>
rect 160 516 202 724
<< poly >>
rect 60 516 202 724
<< ndiff >>
rect 60 516 102 724
<< genericcontact >>
rect -36 -36 276 456
<< genericcontact >>
rect -36 456 276 1076
<< genericcontact >>
rect -94 456 334 1134
<< genericcontact >>
rect -94 -94 334 456
<< genericcontact >>
rect 0 896 240 1040
<< poly >>
rect 0 0 240 144
<< ndiff >>
rect 164 680 204 720
<< pdiff >>
rect 164 680 204 936
<< ndiffusion >>
rect 164 680 204 720
<< pdiffusion >>
rect 164 680 204 720
<< nwell >>
rect 164 680 204 720
<< pwell >>
rect 164 588 204 720
<< via >>
rect 160 104 200 332
<< via >>
rect 160 292 200 350
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 128 416 206 500
<< via >>
rect 44 300 84 640
<< via >>
rect 44 600 110 708
<< metal1 >>
rect 44 300 84 340
<< metal2 >>
rect 44 300 84 340
<< metal3 >>
rect 66 300 106 340
<< metal1 >>
rect 44 300 112 340
<< metal1 >>
rect 48 300 106 340
<< genericcontact >>
rect 0 0 240 1040
<< genericcontact >>
rect 0 896 240 1040
<< poly >>
rect 0 0 240 144
<< ndiff >>
rect 48 300 106 340
<< pdiff >>
rect 44 300 112 340
<< ndiffusion >>
rect 66 300 106 340
<< pdiffusion >>
rect 44 300 84 340
<< nwell >>
rect 44 300 84 340
<< pwell >>
rect 44 600 110 708
<< via >>
rect 44 300 84 640
<< via >>
rect 128 416 206 500
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 160 104 200 144
<< via >>
rect 160 292 200 350
<< via >>
rect 160 104 200 332
<< via >>
rect 164 588 204 720
<< metal1 >>
rect 164 680 204 720
<< metal2 >>
rect 164 680 204 720
<< metal3 >>
rect 164 680 204 720
<< metal1 >>
rect 164 680 204 936
<< metal1 >>
rect 164 680 204 720
<< metal1 >>
rect 140 460 180 500
<< metal1 >>
rect 60 300 100 340
<< end >>