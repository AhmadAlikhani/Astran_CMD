magic
tech scmos
magscale 1 2
timestamp 1687299986
<< m2contact >>
rect 162 570 196 604
<< m2contact >>
rect 160 340 194 374
<< m2contact >>
rect 140 446 174 480
<< m2contact >>
rect 62 570 96 604
<< m2contact >>
rect 60 340 94 374
<< poly >>
rect 118 464 142 488
<< poly >>
rect 116 464 142 672
<< poly >>
rect 118 438 142 462
<< poly >>
rect 118 438 194 488
<< poly >>
rect 116 412 140 462
<< poly >>
rect 116 438 142 462
<< poly >>
rect 114 278 140 436
<< ndiff >>
rect 144 330 210 384
<< ndiff >>
rect 44 330 210 384
<< ndiff >>
rect 44 330 110 384
<< pdiff >>
rect 158 516 200 620
<< pdiff >>
rect 58 516 200 620
<< pdiff >>
rect 58 516 100 620
<< ndiffusion >>
rect -36 -36 276 456
<< pdiffusion >>
rect -36 456 276 1076
<< nwell >>
rect -94 456 334 1134
<< pwell >>
rect -94 -94 334 456
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 570 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 570 208 610
<< metal1 >>
rect 156 104 196 368
<< metal1 >>
rect 156 328 196 386
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 140 434 220 516
<< metal1 >>
rect 56 392 96 598
<< metal1 >>
rect 56 558 96 616
<< metal1 >>
rect 56 392 96 432
<< metal1 >>
rect 56 392 96 432
<< metal1 >>
rect 60 346 100 408
<< metal1 >>
rect 56 368 100 432
<< metal1 >>
rect 60 328 100 386
<< glass >>
rect 0 0 240 1040
<< metal1 >>
rect 0 896 240 1040
<< metal1 >>
rect 0 0 240 144
<< metal1 >>
rect 60 328 100 386
<< metal1 >>
rect 56 368 100 432
<< metal1 >>
rect 60 346 100 408
<< metal1 >>
rect 56 392 96 432
<< metal1 >>
rect 56 392 96 432
<< metal1 >>
rect 56 558 96 616
<< metal1 >>
rect 56 392 96 598
<< metal1 >>
rect 140 434 220 516
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 104 196 144
<< metal1 >>
rect 156 328 196 386
<< metal1 >>
rect 156 104 196 368
<< metal1 >>
rect 150 570 208 610
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 570 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 150 896 190 936
<< metal1 >>
rect 140 460 180 500
<< metal1 >>
rect 60 380 100 420
<< end >>