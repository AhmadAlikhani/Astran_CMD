magic
tech scmos
timestamp 1686702421
input_layout grid
input_grid_coordinates absolute
output_layout absolute
output_grid_coordinates absolute
grid 0.001 0.001
usestrobe
usestamp
<<
<<<
<<<<
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
rect 0 0 4 8
rect 4 0 6 8
rect 6 3 8 5
rect 4 3 6 5
rect 4 0 8 8
rect 2 1 4 7
rect 0 2 2 6
rect 6 2 8 6
rect 0 0 8 8
rect 1 3 2 5
rect 2 2 3 6
rect 3 1 4 7
rect 4 0 5 8
rect 5 1 6 7
rect 6 2 7 6
rect 7 3 8 5
rect 8 4 9 4
